module top #()
();

  enumt dut ();

endmodule : top
