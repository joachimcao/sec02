module top #()
();

  ter dut ();

endmodule : top
