module top #()
();

  relat dut ();

endmodule : top
