module helloworld (
  // input

  // output

);

  initial begin
    $display("Hello World!");
  end

endmodule : helloworld
