module ter ();


endmodule : ter
