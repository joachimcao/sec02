module top #()
();

  stru dut ();

endmodule : top
