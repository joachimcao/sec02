module top #(
)
(

);

  shifts dut ();

endmodule : top
