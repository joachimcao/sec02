module top #()
();

  conca dut ();

endmodule : top
